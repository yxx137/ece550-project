module mux8to1(A, out);
	input[7:0] A;
	output out;
endmodule